module testbench4;



reg [15:0] x , y , z;
wire [15:0] res1;
wire [15:0] res2;
wire  [127:0] stageX;
wire [127:0] stageY;
wire [127:0] stageZ; 
reg mode;
reg reset = 1;
reg clk = 1'b0;
   
initial
begin
      forever
        #3 clk = !clk;
end


cordic c1( mode, x, y, z, clk, reset, res1, res2, stageX, stageY, stageZ);

initial
begin
	reset = 0;
	#3;
	reset = 1;
end


 
initial begin
	mode <= 0;
     #6
	x <= 16'b0001_1010_0110_0000;  
	y <= 16'b0000_1110_0000_0000;    
	z <= 16'b0000_0010_0000_0000;

	#6
	
	
	x <= 16'b0001_1010_0110_0000;    
	y <= 16'b0000_1110_0000_0000;     
	z <= 16'b1000_0011_0001_0000; 
	
	#6
	
	x <= 16'b1011_1001_1001_0100;    
	y <= 16'b0001_1110_1100_0001;
	z <= 16'b0000_0001_1101_1111;
	 
	#6;
	
	x <= 16'b1011_1001_1001_0100;   
	y <= 16'b0001_1110_1100_0001;  
	z <= 16'b1000_0000_1001_1111;
	 
	#6;
	
	x <= 16'b1000_1010_0010_1101;   
	y <= 16'b1000_1000_0010_0000;		
	z <= 16'b0000_0000_0000_1000;
	
	#6
	
	x <= 16'b1000_1010_0010_1101; 
	y <= 16'b1000_1000_0010_0000;      
	z <= 16'b1000_0010_0100_1000;
	
	#6
	
	x <=  16'b0001_0010_1101_0000;       
	y <=  16'b1001_0000_0000_0000;     
	z <=  16'b1000_0000_1111_1111;
	 
	#6

	x <=  16'b0001_0010_1101_0000;      
	y <=  16'b1001_0000_0000_0000;	   
	z <=  16'b0000_0000_1111_1111;
end  

initial 
$monitor($time, " res1 = %b res2 = %b",  res1 , res2);


endmodule

